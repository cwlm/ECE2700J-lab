module roller

endmodule